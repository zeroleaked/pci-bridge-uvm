`ifndef PCI_BRIDGE_TB_TOP
`define PCI_BRIDGE_TB_TOP
 `include "uvm_macros.svh"
`include "pci_bridge_pci_interface.sv"
import uvm_pkg::*;
module pci_bridge_tb_top;
	 
 
	import pci_bridge_test_list::*;

	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Local Fields
	//////////////////////////////////////////////////////////////////////////////
	parameter cycle = 30 ;
	bit clk;
	//////////////////////////////////////////////////////////////////////////////
	//clock generation
	//////////////////////////////////////////////////////////////////////////////
	initial begin
		 clk=0;
		 forever #(cycle/2) clk=~clk;
	end
	//////////////////////////////////////////////////////////////////////////////
	//creatinng instance of interface, inorder to connect DUT and testcase
	//////////////////////////////////////////////////////////////////////////////
	pci_bridge_pci_interface pci_intf(clk);
	
	//////////////////////////////////////////////////////////////////////////////
	/*********************pci_bridge DUT Instantation **********************************/
	//////////////////////////////////////////////////////////////////////////////


	TOP dut_inst(
		.CLK(clk),
		.AD(pci_intf.AD),
		.CBE(pci_intf.CBE),
		.RST(pci_intf.RST),
		.INTA(pci_intf.INTA),
		.REQ(pci_intf.REQ),
		.GNT(pci_intf.GNT),
		.FRAME(pci_intf.FRAME),
		.IRDY(pci_intf.IRDY),
		.IDSEL(pci_intf.IDSEL),
		.DEVSEL(pci_intf.DEVSEL),
		.TRDY(pci_intf.TRDY),
		.STOP(pci_intf.STOP),
		.PAR(pci_intf.PAR),
		.PERR(pci_intf.PERR),
		.SERR(pci_intf.SERR)
	);


	
	//////////////////////////////////////////////////////////////////////////////
	/*********************starting the execution uvm phases**********************/
	//////////////////////////////////////////////////////////////////////////////
	initial begin
		run_test();
	end
	//////////////////////////////////////////////////////////////////////////////
	/**********Set the Interface instance Using Configuration Database***********/
	//////////////////////////////////////////////////////////////////////////////
	initial begin
		uvm_config_db#(virtual pci_bridge_pci_interface)::set(uvm_root::get(),"*","intf",pci_intf);
	end

endmodule

`endif



