`ifndef WB_WRITE_SEQ
`define WB_WRITE_SEQ
class wb_write_seq extends wb_api_base_seq;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Sequence utils
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(wb_write_seq)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new
	// Description : sequence constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "wb_write_seq");
		super.new(name);
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : set_address 
	// Description : override base set_address 
	//////////////////////////////////////////////////////////////////////////////
	task set_address(input bit [31:0] address);
		this.req_address = address | W_BASE_ADDR_1;
	endtask
	///////////////////////////////////////////////////////////////////////////////
	// Method name : do_randomize 
	// Description : Setup randomize constraints for config read
	//////////////////////////////////////////////////////////////////////////////
	function bit do_randomize();
		return req.randomize() with {
			req.is_write == 1'b1;
			req.address[31:2] == req_address[31:2];
			req.data == req_data;
			req.select == 4'hF;
		};
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : write_transaction
	// Description : do a write wb transaction
	//////////////////////////////////////////////////////////////////////////////
	task write_transaction(input bit [31:0] address, data);
		set_address(address);
		req_data = data;
		is_write = 1;
		start(sequencer);
	endtask
	 
endclass

`endif

