`ifndef PCI_CONFIG_TRANSACTION 
`define PCI_CONFIG_TRANSACTION

class pci_config_transaction extends uvm_sequence_item;
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction fields
	//////////////////////////////////////////////////////////////////////////////
	rand bit [31:0] address;
	rand bit [3:0] command;
	rand bit [31:0] data;
	rand bit is_write;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils_begin(pci_config_transaction)
		`uvm_field_int(address, UVM_ALL_ON)
		`uvm_field_int(command, UVM_ALL_ON)
		`uvm_field_int(data, UVM_ALL_ON)
		`uvm_field_int(is_write, UVM_ALL_ON)
	`uvm_object_utils_end
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_config_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////

	//////////////////////////////////////////////////////////////////////////////
	// Method name : drive_address_phase();
	// Description : PCI drive address phase
	//////////////////////////////////////////////////////////////////////////////
	task drive_address_phase(virtual pci_bridge_pci_interface vif);
		vif.dr_cb.FRAME <= 1'b0;	// Assert FRAME#
		vif.dr_cb.AD <= address;
		vif.dr_cb.CBE <= command;
		vif.dr_cb.IDSEL <= 1'b1;	// Assert IDSEL for config space access
	endtask
	//////////////////////////////////////////////////////////////////////////////
	// Method name : wait_for_target();
	// Description : PCI data phase wait for target ready
	//////////////////////////////////////////////////////////////////////////////
	task wait_for_target(virtual pci_bridge_pci_interface vif);
		wait(!vif.dr_cb.DEVSEL && !vif.dr_cb.TRDY);
	endtask
	//////////////////////////////////////////////////////////////////////////////
	// Method name : drive_data_phase();
	// Description : To be overridden by child classes
	//////////////////////////////////////////////////////////////////////////////
	virtual task drive_data_phase(virtual pci_bridge_pci_interface vif);
	endtask
endclass

`endif