`ifndef PCI_BRIGE_WB_TRANSACTION 
`define PCI_BRIGE_WB_TRANSACTION

class wb_transaction extends uvm_sequence_item;
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction fields
	//////////////////////////////////////////////////////////////////////////////
	rand bit is_write;
	rand bit [31:0] address;
	rand bit [31:0] data;
	rand bit [3:0] select;
	rand int trans_id;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils_begin(wb_transaction)
		`uvm_field_int(is_write, UVM_ALL_ON)
		`uvm_field_int(address, UVM_ALL_ON)
		`uvm_field_int(data, UVM_ALL_ON)
		`uvm_field_int(select, UVM_ALL_ON)
		`uvm_field_int(trans_id, UVM_DEFAULT | UVM_NOCOMPARE)
	`uvm_object_utils_end
	 
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "wb_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////
	 
endclass


`endif


