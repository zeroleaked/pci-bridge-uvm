`ifndef PCI_BRIGE_WB_TRANSACTION 
`define PCI_BRIGE_WB_TRANSACTION

class pci_bridge_wb_transaction extends uvm_sequence_item;
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction fields
	//////////////////////////////////////////////////////////////////////////////
	typedef enum {RESET, NORMAL} operation_t;

	operation_t operation;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils_begin(pci_bridge_wb_transaction)
		`uvm_field_enum(operation_t, operation, UVM_ALL_ON)
	`uvm_object_utils_end
	 
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_bridge_wb_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////
	 
endclass


`endif


