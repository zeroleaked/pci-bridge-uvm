`ifndef WB_READ_SEQ
`define WB_READ_SEQ
class wb_read_seq extends wb_api_base_seq;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Sequence utils
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(wb_read_seq)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new
	// Description : sequence constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "wb_read_seq");
		super.new(name);
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : set_address 
	// Description : override base set_address 
	//////////////////////////////////////////////////////////////////////////////
	task set_address(input bit [31:0] address);
		this.req_address = address | W_BASE_ADDR_1;
	endtask
	///////////////////////////////////////////////////////////////////////////////
	// Method name : do_randomize 
	// Description : Setup randomize constraints for config read
	//////////////////////////////////////////////////////////////////////////////
	function bit do_randomize();
		return req.randomize() with {
			req.is_write == 1'b0;
			req.address[31:2] == req_address[31:2];
			req.select == 4'hF;
		};
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : read_transaction
	// Description : do a read wb transaction
	//////////////////////////////////////////////////////////////////////////////
	task read_transaction(input bit [31:0] address);
		set_address(address);
		is_write = 0;
		start(sequencer);
	endtask
	 
endclass

`endif

