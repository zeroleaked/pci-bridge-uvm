`ifndef AGENT_COMMON_PKG
`define AGENT_COMMON_PKG

package agent_common_pkg;
 
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	/////////////////////////////////////////////////////////
	`include "bridge_base_transaction.sv"

endpackage

`endif



