`ifndef PCI_RESPONSE_MEMORY_READ_SEQ
`define PCI_RESPONSE_MEMORY_READ_SEQ
class pci_resp_mem_r_seq extends pci_target_base_seq;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Sequence utils
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(pci_resp_mem_r_seq)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new
	// Description : sequence constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_resp_mem_r_seq");
		super.new(name);
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : do_randomize 
	// Description : Setup randomize constraints for config read
	//////////////////////////////////////////////////////////////////////////////
	function bit do_randomize();
		return req.randomize() with {
			req.data == req_data;
			req.trans_type == PCI_TARGET;
		};
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : read_response
	// Description : do a read pci response
	//////////////////////////////////////////////////////////////////////////////
	task read_response(input bit [31:0] data);
		req_data = data;
		is_write = 0;
		start(sequencer);
	endtask
	 
endclass

`endif


