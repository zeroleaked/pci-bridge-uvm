`ifndef BRIDGE_BASE_TRANSACTION 
`define BRIDGE_BASE_TRANSACTION

class bridge_base_transaction extends uvm_sequence_item;
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction fields
	//////////////////////////////////////////////////////////////////////////////
	// fields for pairing (wb2pci/pci2wb)
	rand bit has_match;
	rand int trans_id;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils_begin(bridge_base_transaction)
		`uvm_field_int(trans_id, UVM_DEFAULT | UVM_NOCOMPARE)
		`uvm_field_int(has_match, UVM_DEFAULT | UVM_NOCOMPARE)
	`uvm_object_utils_end
	 
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "bridge_base_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////
	 
endclass


`endif


