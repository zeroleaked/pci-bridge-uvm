`ifndef PCI_CONFIG_WRITE_TRANSACTION 
`define PCI_CONFIG_WRITE_TRANSACTION

class pci_config_write_transaction extends pci_config_transaction;
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction fields
	//////////////////////////////////////////////////////////////////////////////
	// rand bit [3:0] byte_en;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils_begin(pci_config_write_transaction)
		// `uvm_field_int(byte_en, UVM_ALL_ON)
	`uvm_object_utils_end
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_config_write_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////
	constraint command_c { command == 4'b1011; }
endclass

`endif