`ifndef PCI_BRIDGE_WB_AGENT 
`define PCI_BRIDGE_WB_AGENT

class pci_bridge_wb_agent extends uvm_agent;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of UVC components such as.. driver,monitor,sequencer..etc
	///////////////////////////////////////////////////////////////////////////////
	wb_driver driver;
	wb_sequencer sequencer;
	wb_monitor monitor;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of component utils 
	///////////////////////////////////////////////////////////////////////////////
	`uvm_component_utils(pci_bridge_wb_agent)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new 
	// Description : constructor
	///////////////////////////////////////////////////////////////////////////////
	function new (string name, uvm_component parent);
		super.new(name, parent);
	endfunction : new
	///////////////////////////////////////////////////////////////////////////////
	// Method name : build-phase 
	// Description : construct the components such as.. driver,monitor,sequencer..etc
	///////////////////////////////////////////////////////////////////////////////
	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		driver = wb_driver::type_id::create("driver", this);
		sequencer = wb_sequencer::type_id::create("sequencer", this);
		monitor = wb_monitor::type_id::create("monitor", this);
	endfunction : build_phase
	///////////////////////////////////////////////////////////////////////////////
	// Method name : connect_phase 
	// Description : connect tlm ports ande exports (ex: analysis port/exports) 
	///////////////////////////////////////////////////////////////////////////////
	function void connect_phase(uvm_phase phase);
		driver.seq_item_port.connect(sequencer.seq_item_export);
	endfunction : connect_phase
 
endclass : pci_bridge_wb_agent

`endif
