`ifndef PCI_RESPONSE_MEMORY_READ_SEQ
`define PCI_RESPONSE_MEMORY_READ_SEQ
class pci_resp_mem_r_seq extends pci_target_base_seq;
	bit is_data;
	bit [31:0] req_data;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Sequence utils
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(pci_resp_mem_r_seq)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new
	// Description : sequence constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_resp_mem_r_seq");
		super.new(name);
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : do_randomize 
	// Description : Setup randomize constraints for config read
	//////////////////////////////////////////////////////////////////////////////
	function bit do_randomize();
		return req.randomize() with {
			if (is_data)
				req.data == req_data;
			req.trans_type == PCI_TARGET;
		};
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : read_response
	// Description : do a read pci response
	//////////////////////////////////////////////////////////////////////////////
	task read_response();
		is_write = 0;
		is_data = 0;
		start(sequencer);
	endtask
	///////////////////////////////////////////////////////////////////////////////
	// Method name : read_response_with_data
	// Description : do a read pci response
	//////////////////////////////////////////////////////////////////////////////
	task read_response_with_data(input bit [31:0] data);
		is_write = 0;
		is_data = 1;
		req_data = data;
		start(sequencer);
	endtask
	 
endclass

`endif


