`ifndef BRIDGE_BASE_VSEQ
`define BRIDGE_BASE_VSEQ
class bridge_base_vseq extends uvm_sequence#(uvm_sequence_item);
	uvm_sequencer_base pci_sequencer;
	uvm_sequencer_base wb_sequencer;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Sequence utils
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(bridge_base_vseq)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new
	// Description : sequence constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "bridge_base_vseq");
		super.new(name);
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : body 
	// Description : Body of sequence to send randomized transaction through
	// sequencer to driver
	//////////////////////////////////////////////////////////////////////////////
	virtual task body();
        `uvm_fatal(get_type_name(), "body() not implemented in derived class!")
	endtask
	///////////////////////////////////////////////////////////////////////////////
	// Method name : start_with
	// Description : start with sequencers
	//////////////////////////////////////////////////////////////////////////////
	task start_with(input uvm_sequencer_base pci_sequencer, wb_sequencer);
		this.pci_sequencer = pci_sequencer;
		this.wb_sequencer = wb_sequencer;
		start(null);
	endtask
	 
endclass

`endif


