`ifndef PCI_CONFIG_READ_TRANSACTION 
`define PCI_CONFIG_READ_TRANSACTION

class pci_config_read_transaction extends pci_config_transaction;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(pci_config_read_transaction)
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_config_read_transaction");
		super.new(name);
		is_write = 0;
		command = 4'b1010;	// Config Read command
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Method name : drive_data_phase();
	// Description : PCI data phase of read cycle
	//////////////////////////////////////////////////////////////////////////////
	task drive_data_phase(virtual pci_bridge_pci_interface vif);
		vif.dr_cb.IRDY <= 1'b0;	 // Assert IRDY#
		vif.dr_cb.AD <= 32'bz;		// Release AD bus for target to drive
		vif.dr_cb.CBE <= 4'b0000; // All byte enables active
	endtask
	//////////////////////////////////////////////////////////////////////////////
	// Method name : collect_data();
	// Description : PCI get data from port
	//////////////////////////////////////////////////////////////////////////////
	task collect_data(virtual pci_bridge_pci_interface vif);
		data = vif.dr_cb.AD;
	endtask
endclass

`endif