`ifndef PCI_CONFIG_READ_TRANSACTION 
`define PCI_CONFIG_READ_TRANSACTION

class pci_config_read_transaction extends pci_config_transaction;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(pci_config_read_transaction)
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_config_read_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////
	constraint command_c { command == 4'b1010; }
	constraint is_write_c { is_write == 0; }
endclass

`endif