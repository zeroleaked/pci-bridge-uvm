`ifndef PCI_BRIDGE_WB_MONITOR 
`define PCI_BRIDGE_WB_MONITOR

class pci_bridge_wb_monitor extends uvm_monitor;

	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Virtual interface
	///////////////////////////////////////////////////////////////////////////////
	virtual pci_bridge_wb_interface vif;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Analysis ports and exports 
	///////////////////////////////////////////////////////////////////////////////
	uvm_analysis_port #(pci_bridge_wb_transaction) mon2sb_port;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction item 
	///////////////////////////////////////////////////////////////////////////////
	pci_bridge_wb_transaction act_trans;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of component	utils 
	///////////////////////////////////////////////////////////////////////////////
	`uvm_component_utils(pci_bridge_wb_monitor)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new 
	// Description : constructor
	///////////////////////////////////////////////////////////////////////////////
	function new (string name, uvm_component parent);
		super.new(name, parent);
		act_trans = new();
		mon2sb_port = new("mon2sb_port", this);
	endfunction : new
	///////////////////////////////////////////////////////////////////////////////
	// Method name : build_phase 
	// Description : construct the components
	///////////////////////////////////////////////////////////////////////////////
	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		if(!uvm_config_db#(virtual pci_bridge_wb_interface)::get(this, "", "intf", vif))
			 `uvm_fatal("NOVIF",{"virtual interface must be set for: ",get_full_name(),".vif"});
	endfunction: build_phase
	///////////////////////////////////////////////////////////////////////////////
	// Method name : run_phase 
	// Description : Extract the info from DUT via interface 
	///////////////////////////////////////////////////////////////////////////////
	virtual task run_phase(uvm_phase phase);
		forever begin
			@(vif.rc_cb);
			check_reset_propagation();
			mon2sb_port.write(act_trans);
		end
	endtask : run_phase
	///////////////////////////////////////////////////////////////////////////////
	// Method name : check_reset_propagation
	// Description : Check Wishbone-specific reset conditions
	///////////////////////////////////////////////////////////////////////////////
	bit reset = 0;
	function void check_reset_propagation();
		if (!reset & (vif.rc_cb.RST_O == 1)) begin
			`uvm_info("WB_MONITOR", "Wishbone reset on", UVM_LOW)
			act_trans.operation = pci_bridge_wb_transaction::RESET;
			reset = 1;
		end
		else if (reset & (vif.rc_cb.RST_O == 0)) begin
			`uvm_info("WB_MONITOR", "Wishbone reset off", UVM_LOW)
			act_trans.operation = pci_bridge_wb_transaction::NORMAL;
			reset = 0;
		end
  	endfunction

endclass : pci_bridge_wb_monitor

`endif
