`ifndef PCI_RESPONSE_MEMORY_WRITE_SEQ
`define PCI_RESPONSE_MEMORY_WRITE_SEQ
class pci_resp_mem_w_seq extends pci_target_base_seq;
	///////////////////////////////////////////////////////////////////////////////
	// Declaration of Sequence utils
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils(pci_resp_mem_w_seq)
	///////////////////////////////////////////////////////////////////////////////
	// Method name : new
	// Description : sequence constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_resp_mem_w_seq");
		super.new(name);
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : do_randomize 
	// Description : Setup randomize constraints for config read
	//////////////////////////////////////////////////////////////////////////////
	function bit do_randomize();
		return req.randomize() with {
			req.role == PCI_TARGET;
		};
	endfunction
	///////////////////////////////////////////////////////////////////////////////
	// Method name : write_response
	// Description : do a write pci response
	//////////////////////////////////////////////////////////////////////////////
	task write_response();
		is_write = 1;
		start(sequencer);
	endtask
	 
endclass

`endif


