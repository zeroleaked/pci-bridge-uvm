`ifndef PCI_TRANSACTION 
`define PCI_TRANSACTION

class pci_transaction extends uvm_sequence_item;
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of transaction fields
	//////////////////////////////////////////////////////////////////////////////
	typedef enum bit [3:0] {
		CFG_READ  = 4'b1010,
		CFG_WRITE = 4'b1011,
		MEM_READ  = 4'b0110,
		MEM_WRITE = 4'b0111
	} pci_cmd_t;
	rand pci_cmd_t command;
	rand bit [31:0] address;
	rand bit [31:0] data;
	//////////////////////////////////////////////////////////////////////////////
	//Declaration of Utility and Field macros,
	//////////////////////////////////////////////////////////////////////////////
	`uvm_object_utils_begin(pci_config_transaction)
    	`uvm_field_enum(pci_cmd_t, command, UVM_ALL_ON)
		`uvm_field_int(address, UVM_ALL_ON)
		`uvm_field_int(data, UVM_ALL_ON)
	`uvm_object_utils_end
	//////////////////////////////////////////////////////////////////////////////
	//Constructor
	//////////////////////////////////////////////////////////////////////////////
	function new(string name = "pci_config_transaction");
		super.new(name);
	endfunction
	//////////////////////////////////////////////////////////////////////////////
	// Declaration of Constraints
	//////////////////////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////////
	// Method name : is_write 
	// Description : check if is_write
	///////////////////////////////////////////////////////////////////////////////
	function bit is_write();
		return command[0];
	endfunction
endclass

`endif