`ifndef PCI_BRIDGE_PKG
`define PCI_BRIDGE_PKG

package pci_bridge_pkg;

	`include "pci_bridge_defines.svh" // use this for bench constants

	
endpackage

`endif
