`ifndef PCI_BRIDGE_COVERAGE
`define PCI_BRIDGE_COVERAGE

class pci_bridge_coverage#(type T=pci_bridge_pci_transaction) extends uvm_subscriber#(T);

///////////////////////////////////////////////////////////////////////////////
// Declaration of Local fields
///////////////////////////////////////////////////////////////////////////////
pci_bridge_pci_transaction pci_cov_trans;
`uvm_component_utils(pci_bridge_coverage)
///////////////////////////////////////////////////////////////////////////////
// functional coverage: covergroup for pci
///////////////////////////////////////////////////////////////////////////////
covergroup pci_cg;
	 option.per_instance=1;

	PCI_OPERATION:	coverpoint pci_cov_trans.is_reset { 
					bins reset	= {1};
					bins normal = {0};
				}

endgroup
//////////////////////////////////////////////////////////////////////////////
//constructor
//////////////////////////////////////////////////////////////////////////////
function new(string name="pci_bridge_ref_model", uvm_component parent);
	super.new(name,parent);
	pci_cg =new();
	pci_cov_trans =new();
endfunction
///////////////////////////////////////////////////////////////////////////////
// Method name : sample
// Description : sampling adder_4_bit coverage
///////////////////////////////////////////////////////////////////////////////
function void write(T t);
	this.pci_cov_trans = t;
	pci_cg.sample();
endfunction

endclass

`endif



